library verilog;
use verilog.vl_types.all;
entity gen_circulation is
end gen_circulation;
