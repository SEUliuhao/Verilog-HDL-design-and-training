library verilog;
use verilog.vl_types.all;
entity seg_display_tb is
end seg_display_tb;
