library verilog;
use verilog.vl_types.all;
entity no_block_assign_tb is
end no_block_assign_tb;
