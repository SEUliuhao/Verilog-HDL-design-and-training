library verilog;
use verilog.vl_types.all;
entity data_decrypt_tb is
end data_decrypt_tb;
