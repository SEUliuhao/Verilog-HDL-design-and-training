//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : gate_beh.v
// FUNCTION        : �ŵ�·��ģ��������������ʵ��
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������캽�մ�ѧ������
// UPDATE          :
//******************************************************************************
`timescale 1ns/1ns

module gate_beh
    (
        input i_a, //����5�������ź�
        input i_b,
        input i_c,
        input i_d,
        input i_e,
        
        output o_y //����һ������ź�
    );
    
    //�����ŵ�·֮��������ź�
    reg r_and_o;
    reg r_or1_o;    
    reg r_xor_o;
    reg r_y;
    
    assign o_y = r_y;
    
    
    //��always�����У�����ͼ12-1�ĵ�·�ṹ�������뵽�����˳��
    //��������ֵ�����н�ģ
    
    always @(*) //��ϵ�·��ģ�������ַ�ʽ���������ź��б�������˫�ɱ�����©�����ź�
    begin
        r_and_o = i_a & i_b; //��������ֵ�������Ž��н�ģ
        
        r_or1_o = i_c | i_d; //��������ֵ���Ե�һ�����Ž��н�ģ
        
        r_xor_o = r_and_o ^ r_or1_o; //��������ֵ��������Ž��н�ģ
        
        r_y = r_xor_o | i_e; ////��������ֵ���Եڶ������Ž��н�ģ    
	end
    
endmodule

// END OF gate_beh.v FILE ***************************************************



