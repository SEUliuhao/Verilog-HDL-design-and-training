library verilog;
use verilog.vl_types.all;
entity block_assign_two_tb is
end block_assign_two_tb;
