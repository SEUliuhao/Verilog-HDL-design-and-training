library verilog;
use verilog.vl_types.all;
entity initial_ap is
end initial_ap;
