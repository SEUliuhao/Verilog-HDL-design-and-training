library verilog;
use verilog.vl_types.all;
entity task_gen_clk_app is
end task_gen_clk_app;
