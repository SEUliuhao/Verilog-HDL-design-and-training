library verilog;
use verilog.vl_types.all;
entity gen_special is
end gen_special;
