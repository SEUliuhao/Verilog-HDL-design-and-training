library verilog;
use verilog.vl_types.all;
entity hdb3_code_tb is
end hdb3_code_tb;
