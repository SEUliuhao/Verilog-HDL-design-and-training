//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : data_encrypt.v
// FUNCTION        : ���ݼ���
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս��
// UPDATE          :
//******************************************************************************

module data_encrypt(
    input i_rst_n,
    input i_clk,
    
    input i_data,       //��������
    output o_code);      //���ܺ�ı������

    
    reg [4 : 0] r_shift;
    
    assign o_code = r_shift[4];
    
//*********************************PROCESS**************************************
// FUNCTION        :����ͼ14-1�Ľṹ�������ݼ���
//******************************************************************************     
    always @(negedge i_rst_n, posedge i_clk)
    begin
        if(~i_rst_n)
        begin
            r_shift <= 5'b0;
        end
        else
        begin
            r_shift[3 : 0] <= r_shift[4 : 1];
            r_shift[4] <= r_shift[0] ^ r_shift[2] ^ i_data;
        end
    end
endmodule

// END OF data_encrypt.v FILE *********************************************************
                 
       
            
    
    