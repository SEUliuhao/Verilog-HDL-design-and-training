library verilog;
use verilog.vl_types.all;
entity spi_slave_tb is
end spi_slave_tb;
