library verilog;
use verilog.vl_types.all;
entity timing_block_assign_two_tb is
end timing_block_assign_two_tb;
