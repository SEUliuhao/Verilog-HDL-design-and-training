//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : mux2to1.v
// FUNCTION        : 2ѡ1������
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս��
// UPDATE          :
//******************************************************************************

module mux2to1(
	input A,
	input B,
	input sel,
	
	output reg Y
);

//*********************************always***************************************
// FUNCTION        :����sel��ֵѡ������ź�Y��A����B
//****************************************************************************** 
    always @(A, B, sel)
    begin
        if(sel)
            Y = B;
        else
            Y = A;
    end
endmodule
// END OF mux2to1.v FILE *******************************************************
           