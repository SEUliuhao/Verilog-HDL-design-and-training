library verilog;
use verilog.vl_types.all;
entity display_write_task is
end display_write_task;
