//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : half_adder.v
// FUNCTION        : ��ӷ�����ģ
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������պ����ѧ������
// UPDATE          :
//******************************************************************************
module half_adder(
    input I_a,      //����1
    input I_b,      //����2
    
    output O_sum,   //��
    output O_cout   //��λ�ź�
);


//*********************************PROCESS**************************************
// FUNCTION        :��ӷ������߼�ʵ��
//****************************************************************************** 
    assign O_sum = I_a ^ I_b;
    assign O_cout = I_a & I_b;
    
endmodule


