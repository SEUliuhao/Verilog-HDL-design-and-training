library verilog;
use verilog.vl_types.all;
entity crc_one_tb is
end crc_one_tb;
