
//*******************************FILE HEAD**************************************
//*********************?Verilog HDL ???????????*********************
// FILE NAME       : counter_tbt.v
// FUNCTION        : counter.vģ��Ĳ���ƽ̨
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������պ����ѧ������
// UPDATE					 : 
//******************************************************************************
`timescale 1ns/1ns

module counter_tb();
    
    reg rst_n;
    reg clk;
    
    wire [7 : 0] cnt;
    wire cout;

//ʵ����������ģ��counter    
    counter I1_counter(
        .I_rst_n(rst_n),
        .I_clk(clk),
        .O_cnt(cnt),
        .O_cout(cout)
        );

//*********************************PROCESS**************************************
// FUNCTION        :��ʼ��ʱ���ź�clk����λ�ź�rst_n
//******************************************************************************        
    initial
    begin
        clk = 1'b0;
        rst_n = 1'b0;
        #4 rst_n = 1'b1;
    end
    
//*********************************PROCESS**************************************
// FUNCTION        :��������Ϊ2ns��ʱ���ź�
//******************************************************************************    
    always #1 clk <= ~clk;
    
endmodule
// END OF count.v FILE *********************************************************


        
        