library verilog;
use verilog.vl_types.all;
entity demux1to4_tb is
end demux1to4_tb;
