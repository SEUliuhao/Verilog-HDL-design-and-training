library verilog;
use verilog.vl_types.all;
entity data_encrypt_tb is
end data_encrypt_tb;
