library verilog;
use verilog.vl_types.all;
entity file_input_task is
end file_input_task;
