//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : data_decrypt_tb.v
// FUNCTION        : ���ݽ���ģ�����ƽ̨
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս��
// UPDATE          :
//******************************************************************************
`timescale 1ns/1ns

module data_decrypt_tb();      

    
    reg r_rst_n;
    reg r_clk;
    reg r_data;
    
    wire w_code;    //����������� 
    wire w_data;    //�����������
   
//*********************************PROCESS**************************************
// FUNCTION        :��ʼ��r_rst_n
//******************************************************************************     
    initial
    begin
            r_rst_n = 1'b0;
        #10 r_rst_n = 1'b1; 
    end

//*********************************PROCESS**************************************
// FUNCTION        :��ʼ��r_clk,��������Ϊ2ns��ʱ���ź�
//******************************************************************************     
    initial
    begin
            r_clk = 1'b0;
        forever
            #1  r_clk = ~r_clk;
    end
//*********************************PROCESS**************************************
// FUNCTION        :��ʼ��r_data���������0��1����
//******************************************************************************     
    initial
    begin
            r_data = 1'b0;
        forever
            #2  r_data = $random % 2;
    end

//*********************************PROCESS**************************************
// FUNCTION        :ʵ��������ģ��data_encrypt
//******************************************************************************     
    data_encrypt I1_data_encrypt(
                                    .i_rst_n(r_rst_n),
                                    .i_clk(r_clk),
                                    .i_data(r_data),
                                    .o_code(w_code)
                                 );

//*********************************PROCESS**************************************
// FUNCTION        :ʵ��������ģ��data_encrypt
//******************************************************************************     
    data_decrypt I1_data_decrypt(
                                    .i_rst_n(r_rst_n),
                                    .i_clk(r_clk),
                                    .i_code(w_code),    
                                    .o_data(w_data)
                                 );                                 
                                 
    
endmodule
// END OF data_encrypt.v FILE *********************************************************
                 
       
            
    
    