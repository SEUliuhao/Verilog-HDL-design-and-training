library verilog;
use verilog.vl_types.all;
entity jk_trig_tb is
end jk_trig_tb;
