//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : crc_three_tb.v
// FUNCTION        : CRC���뷽ʽ��ģ�����ƽ̨
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս��
// UPDATE          :
//******************************************************************************
`timescale 1ns/1ns

module crc_three_tb();      
    
    reg [2 : 0] r_data;
    
    wire [3 : 0] w_crc_code;    //CRC�����ź� 

       

//*********************************PROCESS**************************************
// FUNCTION        :��ʼ��r_data
//******************************************************************************     
    initial
    begin
            r_data = 1'b0;
        forever
            #1  r_data = r_data + 3'd1;
    end

//*********************************PROCESS**************************************
// FUNCTION        :ʵ����CRC����ģ��crc_three
//******************************************************************************     
    crc_three I1_crc_three(
                        .i_data(r_data),
                        .o_crc_code(w_crc_code)
                      );
    
endmodule
// END OF data_encrypt.v FILE *********************************************************
                 
       
            
    
    

