library verilog;
use verilog.vl_types.all;
entity file_output_task is
end file_output_task;
