library verilog;
use verilog.vl_types.all;
entity decoder4to10_tb is
end decoder4to10_tb;
