library verilog;
use verilog.vl_types.all;
entity gate_consctruct_tb is
end gate_consctruct_tb;
