library verilog;
use verilog.vl_types.all;
entity gate_dataflow_tb is
end gate_dataflow_tb;
