library verilog;
use verilog.vl_types.all;
entity always_app is
end always_app;
