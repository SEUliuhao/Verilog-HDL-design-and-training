//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : assign_app_two.v
// FUNCTION        : ��ʾӦ��assign������ֵ���ʵ��˫��˿ڵĲ���
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������պ����ѧ������
// UPDATE          :
//******************************************************************************

module assign_app_two(
    input din, //�������룬��˫��˿�д������
    input wr,  //˫��˿ڵĶ�д�����ź�,�͵�ƽΪд���ߵ�ƽΪ��
    
    output dout, //�����������˫��˿ڶ���������
    
    inout data   //˫��˿�
    );
    
//Ӧ��assign������ֵ���ʵ��˫�˿ڵĶ�д����
//��˫�˿�д����
    assign data = (~wr)? din : 1'bz;
//�Ӷ˿ڶ�����
    assign dout = data;
//�Դ�˫��˿ڶ�����������Ҫ����wr�ź�����һЩ�жϡ�
//ֻ����wrΪ�ߵ�ʱ��doutֵ����˫��˿�data��ֵ������doutֵΪdin��ֵ

endmodule
// END OF assign_app_two.v FILE *********************************************************     
