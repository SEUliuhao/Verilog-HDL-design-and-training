library verilog;
use verilog.vl_types.all;
entity arithmetic_op is
end arithmetic_op;
