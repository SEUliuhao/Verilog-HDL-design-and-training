library verilog;
use verilog.vl_types.all;
entity hdb3_decode_tb is
end hdb3_decode_tb;
