library verilog;
use verilog.vl_types.all;
entity task_app is
end task_app;
