//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : gate_dataflow.v
// FUNCTION        : �ŵ�·��ģ��������������ʵ��
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������캽�մ�ѧ������
// UPDATE          :
//******************************************************************************
`timescale 1ns/1ns

module gate_dataflow
    (
        input i_a, //����5�������ź�
        input i_b,
        input i_c,
        input i_d,
        input i_e,
        
        output o_y //����һ������ź�
    );
    
    //�����ŵ�·֮��������ź�
    wire w_and_o;
    wire w_or1_o;    
    wire w_xor_o;
    
    //����ͼ12-1�ĵ�·�ṹ�������뵽�����˳��
    //��������ֵ�����н�ģ
    
    assign w_and_o = i_a & i_b; //��������ֵ�������Ž��н�ģ
    
    assign w_or1_o = i_c | i_d; //��������ֵ���Ե�һ�����Ž��н�ģ
    
    assign w_xor_o = w_and_o ^ w_or1_o; //��������ֵ��������Ž��н�ģ
    
    assign o_y = w_xor_o | i_e; //��������ֵ���Եڶ������Ž��н�ģ 
   
    
endmodule

// END OF gate_dataflow.v FILE ***************************************************



