library verilog;
use verilog.vl_types.all;
entity monitor_task is
end monitor_task;
