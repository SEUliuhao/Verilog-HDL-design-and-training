library verilog;
use verilog.vl_types.all;
entity d_trig_tb is
end d_trig_tb;
