
module noblock_assign
    (
        input a,
        input b, 
        input c,
        input d,
        
        output y
    );
    
    reg y_r;
    reg temp1;
    reg temp2;
    assign y = y_r;
    
    always @(a, b, c, d)
    begin
        temp1 = a & b;
        temp2 = c ^ d;
        y_r = temp1 | temp2;
    end
    
endmodule


