library verilog;
use verilog.vl_types.all;
entity gate_beh_tb is
end gate_beh_tb;
