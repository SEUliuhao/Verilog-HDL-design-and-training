library verilog;
use verilog.vl_types.all;
entity crc_three_tb is
end crc_three_tb;
