//*******************************FILE HEAD**************************************
//*********************��Verilog HDL �����ʵս������Դ����*********************
// FILE NAME       : decoder4to10.v
// FUNCTION        : 4λ���ݵ�10λ���ص�������
// AUTHOR          : 
// DATE & REVISION : 
// COMPANY         : ��Verilog HDL �����ʵս�����������������캽�մ�ѧ������
// UPDATE          :
//******************************************************************************
`timescale 1ns/1ns

module decoder4to10
    (
        input [3: 0]i_data, //����10λ����������        
        
        output [9 : 0] o_decode //����4λ�ı������
    );
    
    //��������ź�o_code�Ļ���
    reg [9 :0] r_decode;
    
    assign o_decode = r_decode; //ͨ��assign������ֵ�����±������
    
       
   
    always @(*) //ʹ��always���̵���Ϊ��ʽ�����ȽϷ���
    begin
   	    case(i_data)
   	        4'b0001: r_decode = 10'b0000000001; //��ϵ�·ʹ��������ֵ���
   	        4'b0010: r_decode = 10'b0000000010;
   	        4'b0011: r_decode = 10'b0000000100;
   	        4'b0100: r_decode = 10'b0000001000;
   	        4'b0101: r_decode = 10'b0000010000;
   	        4'b0110: r_decode = 10'b0000100000;
   	        4'b0111: r_decode = 10'b0001000000;
   	        4'b1000: r_decode = 10'b0010000000;
   	        4'b1001: r_decode = 10'b0100000000;
   	        4'b1010: r_decode = 10'b1000000000;
   	        default: r_decode = 10'b0000000000; //��Ҫ����Ĭ�Ϸ�֧�ĸ�ֵ���������������
   	    endcase
	end
    
endmodule

// END OF decoder4to10.v FILE ***************************************************



