library verilog;
use verilog.vl_types.all;
entity strobe_task is
end strobe_task;
