library verilog;
use verilog.vl_types.all;
entity function_app is
end function_app;
