library verilog;
use verilog.vl_types.all;
entity simulation_time_task is
end simulation_time_task;
