library verilog;
use verilog.vl_types.all;
entity crc_two_tb is
end crc_two_tb;
