library verilog;
use verilog.vl_types.all;
entity noblock_assign_tb is
end noblock_assign_tb;
