library verilog;
use verilog.vl_types.all;
entity printtimescale_task is
end printtimescale_task;
