library verilog;
use verilog.vl_types.all;
entity coder10to4_tb is
end coder10to4_tb;
